`define RESET_PC 32'h00000000
